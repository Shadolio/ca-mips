module register_5 (wordOut, wordIn, write, reset, clk);
	input write, reset, clk;
	input [4:0] wordIn;
	output reg [4:0] wordOut;

	always @(posedge clk, posedge reset) begin

		if(reset) wordOut <= 4'd0;

		else if(write) wordOut <= wordIn;

	end

endmodule

module register_5_tb ();
	reg write, reset, clk;
	reg [4:0] wordIn;
	wire [4:0] wordOut;

	register_5 testReg (wordOut, wordIn, write, reset, clk);

	initial begin

		$monitor("In: %h, Out: %h", wordIn, wordOut);

		#5 reset <= 1;

		#5 wordIn <= 4'd5;

		write <= 1;
		reset <= 0;
		#5 clk <= 1;

	end

endmodule
