module mips_proc ();

	initial begin
		#10 $display("MIPS processor starting...");
		#10 $display("Welcome to MIPS processor!");
	end

endmodule
